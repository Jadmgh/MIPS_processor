library verilog;
use verilog.vl_types.all;
entity test_alucontrol_vlg_vec_tst is
end test_alucontrol_vlg_vec_tst;
