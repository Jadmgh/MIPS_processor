library verilog;
use verilog.vl_types.all;
entity Control_testing_vlg_vec_tst is
end Control_testing_vlg_vec_tst;
