library verilog;
use verilog.vl_types.all;
entity testing_reg_file_vlg_vec_tst is
end testing_reg_file_vlg_vec_tst;
