library verilog;
use verilog.vl_types.all;
entity test_edgedetector_vlg_vec_tst is
end test_edgedetector_vlg_vec_tst;
