library verilog;
use verilog.vl_types.all;
entity test_alucontrol_vlg_check_tst is
    port(
        op              : in     vl_logic_vector(2 downto 0);
        sampler_rx      : in     vl_logic
    );
end test_alucontrol_vlg_check_tst;
