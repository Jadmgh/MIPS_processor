library verilog;
use verilog.vl_types.all;
entity testing_alu_vlg_vec_tst is
end testing_alu_vlg_vec_tst;
